// Code your testbench here
// or browse Examples
`include "palindrome_tb.sv";